----------------------------------------------------------------------------------
-- This Component are made to generate integral image
-- Designer : Jason Danny Setiawan
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ii_gen_top is
	Port ( clk 					: in STD_LOGIC; 								-- Typical 100 MHz clock
			 reset			 	: in STD_LOGIC; 								-- reset
			 ii_start			: in STD_LOGIC; 								-- Generated by top level FSM
			 din					: in STD_LOGIC_VECTOR(11 downto 0); 	-- Data 12 bit image from main buffer
			 image_scale		: in STD_LOGIC_VECTOR(1 downto 0); 		-- Scaling image
			 scaleImg_x_base	: in STD_LOGIC_VECTOR(5 downto 0); 		-- x base position of integral image -> 64 max
			 scaleImg_y_base	: in STD_LOGIC_VECTOR(5 downto 0);		-- y base position of integral image -> 48 max
			 mem_state			: in STD_LOGIC;								-- ii_buffer partition selector
			 ii_data_in			: in STD_LOGIC_VECTOR(18 downto 0);		-- feedback berisi integral image from prev row
			 iix2_data_in		: in STD_LOGIC_VECTOR(22 downto 0);		-- feedback berisi squared integral image from prev row
			 
			 ii_wren				: out STD_LOGIC;								-- buffer write enable
			 ii_address			: out STD_LOGIC_VECTOR (11 downto 0); 	-- address ii dan iix2 buffer
			 
			 ii_data_o			: out STD_LOGIC_VECTOR(18 downto 0);	-- data output to ii buffer
			 iix2_data_o		: out STD_LOGIC_VECTOR(22 downto 0);	-- data output to iix2 buffer
			 image_rdaddress	: out STD_LOGIC_VECTOR(13 downto 0);	-- address for requesting data from main buffer
			 done					: out STD_LOGIC);
end ii_gen_top;

architecture Behavioral of ii_gen_top is

component rgb2grey
	Port ( Datain : in  STD_LOGIC_VECTOR (11 downto 0);
          Dataout : out  STD_LOGIC_VECTOR (7 downto 0));
end component rgb2grey;

constant II_WIDTH : unsigned(5 downto 0) := to_unsigned(50,6);
constant II_HEIGHT : unsigned(5 downto 0) := to_unsigned(40,6);

-- x pos relative to ii ( 0 - 49 )
signal x : std_logic_vector(5 downto 0);
signal x_count_reset : std_logic;
signal x_count_en : std_logic;

-- y pos relative to ii ( 0 - 39 )
signal y : std_logic_vector(5 downto 0);
signal y_count_reset : std_logic;
signal y_count_en : std_logic;

-- scaled image address
signal image_address_base : std_logic_vector (13 downto 0) := (others => '0');

-- image rd address
signal address_accu_reset : std_logic := '0';
signal image_rdaddress_reg : std_logic_vector(13 downto 0):=(others=>'0');
signal image_address_base_reg : std_logic_vector(13 downto 0):=(others=>'0');
-- gray data declaration
signal gray_data : std_logic_vector(7 downto 0);
signal gray_data_square : std_logic_vector(15 downto 0);
signal gray_data_square_per16 : std_logic_vector(11 downto 0);

-- mini state machine:
---- since the last scale is 41.67%, the image must be resize to its 12/5 original size
---- that means I should sample 5 pixel, from original 12 pixels.
------- If I use simple addition by 2 (skip a pixel after another) there will be 6 pixel sampled
------- out of 12. That is 50% resizing. Same thing happens in addition by 3 and make 33% resizing.
----	I need to add by 1 and by 2 respectively, so i need these state to sample with that method.

type state_parity is (odd, even);
signal state_oddeven : state_parity := odd;
signal state_oddeveny : state_parity := odd;


signal addr_base_temp1 : std_logic_vector (13 downto 0);
signal addr_base_temp2 : std_logic_vector (13 downto 0); 

-- These value needs to be added to original image address
-- So, if I scan x*y pixels, then after x pixel i should move to the max_x+1 pixels and so on,
--	then i need a value to jump from x to max_x + 1
-- Formula : (max_img_width - ii_width - 1)*scale
-- II dimension : 50 x 40 = 2000
type lut is array ( 0 to 3 ) of std_logic_vector(8 downto 0);
constant my_lut : lut := ( std_logic_vector(to_unsigned(0, 9)), -- not used
                           std_logic_vector(to_unsigned(256, 9)),  -- (128 - 50 - 1) * 2 = 154
                           std_logic_vector(to_unsigned(384, 9)),  -- (128 - 50 - 1) * 3 = 231
									std_logic_vector(to_unsigned(0, 9)));  
signal arrival : std_logic_vector(8 downto 0); -- output signal of my_lut0 process

signal ii_wraddress : std_logic_vector(11 downto 0);
signal ii_rdaddress : std_logic_vector(11 downto 0);

signal ii_address_sel  : std_logic;

signal xbase_ori_1  	: std_logic_vector(6 downto 0);
signal xbase_ori_2 	: std_logic_vector(11 downto 0);
signal xbase_ori_2a 	: std_logic_vector(11 downto 0);
signal xbase_ori_2b 	: std_logic_vector(11 downto 0);
signal xbase_ori_2c 	: std_logic_vector(11 downto 0);
signal xbase_ori_2d 	: std_logic_vector(11 downto 0);
signal xbase_ori	 	: std_logic_vector(6 downto 0);
signal ybase_ori_1 	: std_logic_vector(6 downto 0);
signal ybase_ori_2 	: std_logic_vector(11 downto 0);
signal ybase_ori_2a	: std_logic_vector(11 downto 0);
signal ybase_ori_2b	: std_logic_vector(11 downto 0);
signal ybase_ori_2c	: std_logic_vector(11 downto 0);
signal ybase_ori_2d	: std_logic_vector(11 downto 0);
signal ybase_ori	 	: std_logic_vector(6 downto 0);

signal sum : std_logic_vector(13 downto 0);
signal sum2 : std_logic_vector(17 downto 0);
signal sum_extend : std_logic_vector(18 downto 0);
signal sum2_extend : std_logic_vector(22 downto 0);
signal sum3 : std_logic_vector(18 downto 0);
signal sum4 : std_logic_vector(22 downto 0);

signal ii_data_accu : std_logic_vector(13 downto 0); -- accumulator register out
signal iix2_data_accu : std_logic_vector(17 downto 0); -- accumulator register out (squared)

signal ii_data_o_s : std_logic_vector(18 downto 0);
signal iix2_data_o_s : std_logic_vector(22 downto 0);

-- Temporary Register
-- Register 0
signal reg0_x : std_logic_vector(5 downto 0);
signal reg0_y : std_logic_vector(5 downto 0);
signal reg0_ii_wraddress : std_logic_vector(11 downto 0);
signal reg0_image_data : std_logic_vector(11 downto 0);
signal reg0_ii_data : std_logic_vector(18 downto 0);
signal reg0_iix2_data : std_logic_vector(22 downto 0);
signal reg0_accu_reset : std_logic;
signal reg0_accu_en : std_logic;
signal reg0_done : std_logic;

-- Register 1
signal reg1_x : std_logic_vector(5 downto 0);
signal reg1_y : std_logic_vector(5 downto 0);
signal reg1_ii_wraddress : std_logic_vector(11 downto 0);
signal reg1_gray_data : std_logic_vector(7 downto 0);
signal reg1_ii_data : std_logic_vector(18 downto 0);
signal reg1_iix2_data : std_logic_vector(22 downto 0);
signal reg1_accu_reset : std_logic;
signal reg1_accu_en : std_logic;
signal reg1_done : std_logic;

-- R2
signal reg2_x : std_logic_vector(5 downto 0);
signal reg2_y : std_logic_vector(5 downto 0);
signal reg2_ii_wraddress : std_logic_vector(11 downto 0);
signal reg2_gray_data : std_logic_vector(7 downto 0);
signal reg2_gray_data_square : std_logic_vector(11 downto 0);
signal reg2_ii_data : std_logic_vector(18 downto 0);
signal reg2_iix2_data : std_logic_vector(22 downto 0);
signal reg2_accu_reset : std_logic;
signal reg2_accu_en : std_logic;
signal reg2_done : std_logic;

-- R3
signal reg3_x : std_logic_vector(5 downto 0);
signal reg3_y : std_logic_vector(5 downto 0);
signal reg3_ii_wraddress : std_logic_vector(11 downto 0);
signal reg3_sum_extend : std_logic_vector(18 downto 0);
signal reg3_sum2_extend : std_logic_vector(22 downto 0);
signal reg3_sum3 : std_logic_vector(18 downto 0);
signal reg3_sum4 : std_logic_vector(22 downto 0);
signal reg3_done : std_logic;
  
signal reset_done_reg : std_logic;
signal done_reg : std_logic;

signal accu_reset : std_logic;
signal accu_en : std_logic;

signal pipeline_step : std_logic;
signal pipeline_reset	: std_logic;

type STATE_TYPE is (state_RESET, latch_RAM_read, latch_RAM_write, SOFT_reset, state_DONE);
signal state,next_state : STATE_TYPE;

signal buffer_write_en : std_logic;
signal done_s : std_logic;

begin
rgb2grey_inst : rgb2grey port map (
	Datain => reg0_image_data,
	Dataout => gray_data);
	
gray_data_square <= std_logic_vector(unsigned(reg1_gray_data)*unsigned(reg1_gray_data));
gray_data_square_per16 <= gray_data_square(15 downto 4);

x_counter : process (clk, x_count_reset, x_count_en) begin
	if (x_count_reset = '1')then
		x <= (others => '0');
	elsif (rising_edge(clk) and (x_count_en = '1')) then
		x <= std_logic_vector(unsigned(x)+to_unsigned(1,6));
	end if;
end process x_counter;
	
y_counter : process (clk, y_count_reset, y_count_en) begin
	if (y_count_reset = '1')then
		y <= (others => '0');
	elsif (rising_edge(clk) and (y_count_en = '1')) then
		y <= std_logic_vector(unsigned(y)+to_unsigned(1,6));
	end if;
end process y_counter;

-- Calculate the position of integral image in original 128x96 image.
-- Scaling used : 50% 41.67% 
xbase_ori_1 <= scaleImg_x_base & '0';

xbase_ori_2a <= scaleImg_x_base & "000000";
xbase_ori_2b <= "000" & scaleImg_x_base & "000";
xbase_ori_2c <= "0000" & scaleImg_x_base & "00";
xbase_ori_2d <= "000000" & scaleImg_x_base;
xbase_ori_2 <= std_logic_vector(unsigned(xbase_ori_2a) + unsigned(xbase_ori_2b) + unsigned(xbase_ori_2c) + unsigned(xbase_ori_2d));

ybase_ori_1 <= scaleImg_y_base & '0';

ybase_ori_2a <= scaleImg_y_base & "000000";
ybase_ori_2b <= "000" & scaleImg_y_base & "000";
ybase_ori_2c <= "0000" & scaleImg_y_base & "00";
ybase_ori_2d <= "000000" & scaleImg_y_base;
ybase_ori_2 <= std_logic_vector(unsigned(ybase_ori_2a) + unsigned(ybase_ori_2b) + unsigned(ybase_ori_2c) + unsigned(ybase_ori_2d));

process (image_scale,xbase_ori_1,ybase_ori_1,xbase_ori_2,ybase_ori_2) begin
	case (image_scale) is
		when "01" =>
			xbase_ori <= xbase_ori_1(6 downto 0);
			ybase_ori <= ybase_ori_1(6 downto 0);
		
		when "10" =>
			xbase_ori <= xbase_ori_2(11 downto 5);
			ybase_ori <= ybase_ori_2(11 downto 5);
		
		when others =>
			xbase_ori <= (others => '0');
			ybase_ori <= (others => '0');
	end case;
end process;

-- Calculate the position of integral image in scaled image.
-- address base = 128*y + x , 128 is the max pixel in a y (row).
-- Since multipliying 3 digits decimal with 2-3 digits decimal
-- 	take a lot of multipliers. I use this trick
--		address base = 128*y+x
--		128 y = y << 7
--		y = y_ori * scale
--		x = x_ori * scale
addr_base_temp1 <= ybase_ori & "0000000";	-- 7 bit & 7 bit ( *128)
addr_base_temp2 <= "0000000" & xbase_ori; -- 7 bit & 8 bit
image_address_base <= std_logic_vector(unsigned(addr_base_temp1) + unsigned(addr_base_temp2));		
						
arrival <= my_lut(to_integer(unsigned(image_scale)));		

-- image_rdaddress accumulator 
-- (1) since the integral image scans the oringal image, image_address_base specifies the location of the integral image relative to oringal image with scaling adjustments
-- (2) increment the image_rdaddress in a linear scaling fashion 
--     by x_scaled+=image_scale
--     or x_scaled=0, y_scaled+=image_scale											
accu_image_rdaddress: process (clk, address_accu_reset, x_count_en, y_count_en, image_scale, arrival, image_address_base)
  begin
    if rising_edge(clk) then
		if address_accu_reset='1' then
			image_rdaddress_reg <= image_address_base;
			image_address_base_reg <= image_address_base;
		elsif x_count_en='1' then -- address += scale
			if unsigned(image_scale) = 1 then
				image_rdaddress_reg <= std_logic_vector(unsigned(image_rdaddress_reg) + to_unsigned(2,2));
				
			elsif unsigned(image_scale) = 2 then 
				case state_oddeven is
					when even =>
						image_rdaddress_reg <= std_logic_vector(unsigned(image_rdaddress_reg) + unsigned(to_unsigned(3,2)));
						state_oddeven <= odd;
					when odd =>
						image_rdaddress_reg <= std_logic_vector(unsigned(image_rdaddress_reg) + unsigned(to_unsigned(2,2)));
						state_oddeven <= even;
				end case;
			else	
				image_rdaddress_reg <= (others => '0');
			end if;
	 elsif y_count_en='1' then -- address += max_img_width*scale-(ii_width-1)*scale
      if unsigned(image_scale) = 1 then
			image_rdaddress_reg <= std_logic_vector(unsigned(image_address_base_reg) + unsigned(arrival));
			image_address_base_reg <= std_logic_vector(unsigned(image_address_base_reg) + unsigned(arrival));
		
		elsif unsigned(image_scale) = 2 then
			case state_oddeveny is
				when even =>
					image_rdaddress_reg <= std_logic_vector(unsigned(image_address_base_reg) + unsigned(arrival));
					image_address_base_reg <= std_logic_vector(unsigned(image_address_base_reg) + unsigned(arrival));
					state_oddeveny <= odd;
				when odd  =>
					image_rdaddress_reg <= std_logic_vector(unsigned(image_address_base_reg) + to_unsigned(256,8));
					image_address_base_reg <= std_logic_vector(unsigned(image_address_base_reg) + to_unsigned(256,8));
					state_oddeveny <= even;
			end case;
		end if;
    end if;
	end if;
  end process;
  image_rdaddress <= image_rdaddress_reg;
  
  
accu_image_wraddress : process(clk, address_accu_reset, x_count_en, y_count_en) begin
	if rising_edge(clk) then
		if	address_accu_reset='1' then
			if mem_state <= '0' then -- store in upper partition (lower mem)
				ii_wraddress <= (others=>'0');
			else 
				ii_wraddress <= std_logic_vector(to_unsigned(2048,12));
			end if;
		elsif (x_count_en='1' or y_count_en='1') then
			ii_wraddress <= std_logic_vector(unsigned(ii_wraddress) + to_unsigned(1,8));
		end if;
	end if;
end process;
		
-- ii_rdaddress is always ii_mem[x,y-1] = ii_wraddress - II_WIDTH, read previous column value
ii_rdaddress <= std_logic_vector(unsigned(ii_wraddress) - II_WIDTH);
  
-- integral image read and write address share the same buffer address input
address_mux: process (reg3_ii_wraddress, ii_rdaddress, ii_address_sel) begin
	if ii_address_sel='0' then
		ii_address <= ii_rdaddress;
	else
		ii_address <= reg3_ii_wraddress;
	end if;
end process;	

-- accumulator data path
-- gray_data + ii_mem[x,y-1]
sum <= std_logic_vector(unsigned(reg2_gray_data)+unsigned(ii_data_accu)); -- max = 50*255 = 12,750 = 14bit uns 
-- gray_data_square + iix2_mem[x,y-1]
sum2 <= std_logic_vector(unsigned(reg2_gray_data_square)+unsigned(iix2_data_accu)); -- max = 50*4096 = 200,800 = 18bit uns
sum_extend(18 downto 14) <= (others=>'0');
sum_extend(13 downto 0) <= sum;
sum2_extend(22 downto 18) <= (others=>'0');
sum2_extend(17 downto 0) <= sum2;

-- accuulate the ii and iix2 values for a single row at a time
accu_reg: process(clk, reset, reg2_accu_reset, reg2_accu_en, sum, sum2, pipeline_step) begin
	if rising_edge(clk) then
		if (reg2_accu_reset = '1'and pipeline_step = '1') then
			ii_data_accu <= (others=>'0'); -- sync register reset
			iix2_data_accu <= (others=>'0');
		elsif (reg2_accu_en='1' and pipeline_step='1') then -- only accumulate when new data is shifted in pipeline
			ii_data_accu <= sum; -- latch register
			iix2_data_accu <= sum2;
		end if;
	end if;
end process;

sum3 <= std_logic_vector(unsigned(reg2_ii_data)+unsigned(sum));   -- ii_accu + gray_data + ii_mem[x,y-1] 
sum4 <= std_logic_vector(unsigned(reg2_iix2_data)+unsigned(sum2)); -- iix2_accu + gray_data_square + iix2_mem[x,y-1]

-- data output mux .. sel='1' when y=0(dec)
mux0: process(reg3_y,reg3_sum_extend,reg3_sum2_extend,reg3_sum3,reg3_sum4)
begin
	if (reg3_y="000000") then
		ii_data_o_s <= reg3_sum_extend;   -- ii_mem[x,y] <= ii_accu + gray_data
		iix2_data_o_s <= reg3_sum2_extend; -- iix2_mem[x,y] <= iix2_accu + gray_data_square
	else
		ii_data_o_s <= reg3_sum3;   -- ii_mem[x,y] <= ii_accu + gray_data + ii_mem[x,y-1]
		iix2_data_o_s <= reg3_sum4; -- iix2_mem[x,y] <= iix2_accu + gray_data_square + iix2_mem[x,y-1]
   end if;
end process;

-- Pipeline can be used by storing data carried by an integral image (49 x 39) through temporary register
pipeline_process : process (clk, pipeline_reset, pipeline_step, x, y, ii_wraddress, 
									Din, ii_data_in, iix2_data_in, gray_data, gray_data_square,
									sum_extend, sum2_extend, sum3, sum4, accu_reset, accu_en, done_s) begin

	if pipeline_reset = '1' then
		reg0_x				<= (others=>'0');
		reg0_y 				<= (others=>'0');
		reg0_ii_wraddress <= (others=>'0');
		reg0_image_data 	<= (others => '0');
		reg0_ii_data 		<= (others => '0');
		reg0_iix2_data 	<= (others => '0');
		reg0_accu_reset 	<= '1';
		reg0_accu_en 		<= '0';
		reg0_done 			<= '0';
		
		reg1_x 				<= (others => '0');
		reg1_y 				<= (others => '0');
		reg1_ii_wraddress <= (others => '0');
		reg1_gray_data 	<= (others => '0');
		reg1_ii_data 		<= (others => '0');
		reg1_iix2_data 	<= (others => '0');
		reg1_accu_reset 	<= '1';
		reg1_accu_en 		<= '0';
		reg1_done 			<= '0';

		reg2_x 						<= (others => '0');
		reg2_y 						<= (others => '0');
		reg2_ii_wraddress 		<= (others => '0');
		reg2_gray_data 			<= (others => '0');
		reg2_gray_data_square 	<= (others => '0');
		reg2_ii_data 				<= (others => '0');
		reg2_iix2_data 			<= (others => '0');
		reg2_accu_reset 			<= '1';
		reg2_accu_en 				<= '0';
		reg2_done 					<= '0';
		
		reg3_x            <= (others=>'0');
		reg3_y            <= (others=>'0'); 
      reg3_ii_wraddress	<= (others=>'0'); 
      reg3_sum_extend	<= (others=>'0');
      reg3_sum2_extend  <= (others=>'0');
      reg3_sum3         <= (others=>'0');
      reg3_sum4         <= (others=>'0');
      reg3_done         <= '0';
	elsif rising_edge(clk) and pipeline_step = '1' then
		reg0_x				<= x;
		reg0_y 				<= y;
		reg0_ii_wraddress <= ii_wraddress;
		reg0_image_data 	<= Din;
		reg0_ii_data 		<= ii_data_in;
		reg0_iix2_data 	<= iix2_data_in;
		reg0_accu_reset 	<= accu_reset;
		reg0_accu_en 		<= accu_en;
		reg0_done 			<= done_s;
		
		reg1_x 				<= reg0_x;
		reg1_y 				<= reg0_y;
		reg1_ii_wraddress <= reg0_ii_wraddress;
		reg1_gray_data 	<= gray_data;
		reg1_ii_data 		<= reg0_ii_data;
		reg1_iix2_data 	<= reg0_iix2_data;
		reg1_accu_reset 	<= reg0_accu_reset;
		reg1_accu_en 		<= reg0_accu_en;
		reg1_done 			<= reg0_done;

		reg2_x 						<= reg1_x;
		reg2_y 						<= reg1_y;
		reg2_ii_wraddress 		<= reg1_ii_wraddress;
		reg2_gray_data 			<= reg1_gray_data;
		reg2_gray_data_square 	<= gray_data_square_per16;
		reg2_ii_data 				<= reg1_ii_data;
		reg2_iix2_data 			<= reg1_iix2_data;
		reg2_accu_reset 			<= reg1_accu_reset;
		reg2_accu_en 				<= reg1_accu_en;
		reg2_done 					<= reg1_done;
		
		reg3_x            <= reg2_x;
		reg3_y            <= reg2_y; 
      reg3_ii_wraddress	<= reg2_ii_wraddress; 
      reg3_sum_extend	<= sum_extend;
      reg3_sum2_extend  <= sum2_extend;
      reg3_sum3         <= sum3;
      reg3_sum4         <= sum4;
      reg3_done         <= reg2_done;	
	end if;
end process pipeline_process;

statemachine_ctrllr : process (clk, reset, next_state) begin
	if (reset = '1') then
		state <= state_RESET;
	elsif rising_edge(clk) then
		state <= next_state;
	end if;
end process statemachine_ctrllr;

fsm_proc : process (state, ii_start, x, y, ii_address_sel, done_reg) begin
	accu_reset <= '0';
   buffer_write_en <= '0';
   accu_en <= '0';
   x_count_reset <= '0';
   x_count_en <= '0';
   y_count_reset <= '0';
   y_count_en <= '0';
   done_s <= '0';
   ii_address_sel <= '0';
   address_accu_reset <= '0';
   pipeline_step <= '0';
   pipeline_reset <= '0';
   reset_done_reg <= '0';
	
	case state is
		when state_RESET =>
			accu_reset <= '1';
			address_accu_reset <= '1';
			x_count_reset <= '1';
			y_count_reset <= '1';
			pipeline_reset <= '1';
			reset_done_reg <= '1';
			if ii_start = '1' then
				next_state <= latch_RAM_read;
			else
				next_state <= state_RESET;
			end if;
		
		when latch_RAM_read =>
			ii_address_sel <= '0'; --  if ii_address_sel='0' then ii_address <= ii_rdaddress
			next_state <= latch_RAM_write;
		
		when latch_RAM_write =>
			pipeline_step <= '1'; --pipelining active
			buffer_write_en <= '1';
			ii_address_sel <= '1'; -- if ii_address_sel='1' then ii_address <= reg3_iiwrd_addr
		
			if (unsigned(x) = II_WIDTH - to_unsigned(1,6))  then -- ii row accu selesai
				accu_reset <= '1';
				if (unsigned(y) = II_HEIGHT - to_unsigned(1,6)) then -- ii row x line accu selesai
					-- go to done state
						done_s <= '1'; -- flag last pipeline execution with done
						next_state <= state_DONE;
				else
				y_count_en <= '1'; --increment to next ii row
            next_state <= SOFT_reset;
          end if;
        else
          accu_en <= '1'; -- continue to accumulate row ii values
          x_count_en <= '1';
          next_state <= latch_RAM_read;
        end if;
        
      when SOFT_reset =>
        x_count_reset <= '1'; -- sync reset ii x position
        next_state <= latch_RAM_read;
        
      when state_DONE =>
        -- continue to write ii values to buffer unitl done assertion is recieved from last pipeline operation
        if done_reg='1' then
        -- null, stop writing to ii buffer
        else
          ii_address_sel <= '1'; -- setup wraddress
          pipeline_step <= '1'; -- advance remaining pipeline data
          buffer_write_en <= '1';
        end if;
        next_state <= state_DONE; -- stay here, reset at top level
    end case;
  end process;

done_register: process(clk, reset_done_reg, reg3_done)
begin
	if reset_done_reg='1' then
		done_reg <= '0';
	elsif rising_edge(clk) and reg3_done='1' then
		done_reg <= '1';
	end if;
end process;

ii_wren <= buffer_write_en;
ii_data_o <= ii_data_o_s;
iix2_data_o <= iix2_data_o_s;
done <= done_reg;  

end Behavioral;

